`ifndef ALU_PARAMETERS_DEFINE
`define ALU_PARAMETERS_DEFINE

`define ALU_REG_WIDTH 4
`define ALU_USE_PIPELINED_ALPU 0

`endif
