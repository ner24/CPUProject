
module eu_iconIQueue #(
  parameter NUM_CHANNELS = 2,

  //NOTE: in this config, total iqueue size would be IQUEUE_LENGTH * NUM_CHANNELS
  parameter IQUEUE_LENGTH = 4
) (

);


endmodule
