`define VERIF_MODULE_SUFFIX_CONST _simv
`ifdef MODE_SIMULATION
`define MODE_SIM 1
`define VERIF_MODULE_SUFFIX `VERIF_MODULE_SUFFIX_CONST
`else
`define MODE_SIM 0
`define VERIF_MODULE_SUFFIX
`endif

`define SIM_TB_MODULE(m) ``m```VERIF_MODULE_SUFFIX
