module eu_iconIntf import exec_unit_dtypes::*; #(
  
) (
  input  wire type_icon_channel    rx,
  output wire type_icon_rx_channel rx_tx,
  
  output wire type_icon_channel    tx,
  input  wire type_icon_rx_channel tx_rx

  
);



endmodule
