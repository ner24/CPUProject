module eu_iconChannel #(
  parameter NUM_ELEMENTS = 3
) (
  //input wire 
);


endmodule
