module exec_block #(

) (

);


endmodule
