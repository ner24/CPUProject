module Icon_TXQ import exec_unit_dtypes::*; #(

) (
  input  wire clk,
  input  wire reset_n
);

  

endmodule
