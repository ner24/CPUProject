module execution_unit #(

) (

);


endmodule
