module eu_prepop #(

) (

);

  

endmodule
