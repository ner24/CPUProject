`ifndef ALU_PARAMETERS_DEFINE
`define ALU_PARAMETERS_DEFINE

`define ALU_REG_WIDTH 4
`define ALU_USE_PIPELINED_ALPU 0

`define NUM_EXEC_UNITS 2
`define NUM_REG 8

`endif
