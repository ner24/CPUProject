`include "simulation_parameters.sv"
`include "alu_parameters.sv"
