
module eu_iconIQueue import exec_unit_dtypes::*; #(
  parameter NUM_CHANNELS = 2,

  //NOTE: in this config, total iqueue size would be IQUEUE_LENGTH * NUM_CHANNELS
  parameter IQUEUE_LENGTH = 4
) (

);


endmodule
