module alu_front_end #(
  parameter REG_WIDTH = 8
)(
    
);

  

endmodule
