module eu_iconIntf import exec_unit_dtypes::*; #(
  
) (
  inout wire type_icon_channel channel_port
);

  

endmodule
